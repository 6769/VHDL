library verilog;
use verilog.vl_types.all;
entity lab50_vlg_vec_tst is
end lab50_vlg_vec_tst;
