library verilog;
use verilog.vl_types.all;
entity NbitCounter_vlg_vec_tst is
end NbitCounter_vlg_vec_tst;
