library verilog;
use verilog.vl_types.all;
entity multiplexers_vlg_vec_tst is
end multiplexers_vlg_vec_tst;
