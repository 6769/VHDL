library verilog;
use verilog.vl_types.all;
entity Addsub_vlg_vec_tst is
end Addsub_vlg_vec_tst;
