library verilog;
use verilog.vl_types.all;
entity light_vlg_vec_tst is
end light_vlg_vec_tst;
