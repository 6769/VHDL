library verilog;
use verilog.vl_types.all;
entity rotate_shift_register_vlg_vec_tst is
end rotate_shift_register_vlg_vec_tst;
