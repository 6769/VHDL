library verilog;
use verilog.vl_types.all;
entity DiceGame_controller_vlg_vec_tst is
end DiceGame_controller_vlg_vec_tst;
