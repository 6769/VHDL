--
	