library verilog;
use verilog.vl_types.all;
entity light_vlg_check_tst is
    port(
        f               : in     vl_logic;
        g               : in     vl_logic;
        h               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end light_vlg_check_tst;
