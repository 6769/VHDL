library verilog;
use verilog.vl_types.all;
entity View2_vlg_vec_tst is
end View2_vlg_vec_tst;
