library verilog;
use verilog.vl_types.all;
entity counter741_vlg_vec_tst is
end counter741_vlg_vec_tst;
