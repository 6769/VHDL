library verilog;
use verilog.vl_types.all;
entity Control_unit_vlg_vec_tst is
end Control_unit_vlg_vec_tst;
