library verilog;
use verilog.vl_types.all;
entity counter_max10_vlg_vec_tst is
end counter_max10_vlg_vec_tst;
