library verilog;
use verilog.vl_types.all;
entity Game_vlg_vec_tst is
end Game_vlg_vec_tst;
