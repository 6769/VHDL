library verilog;
use verilog.vl_types.all;
entity View_output_vlg_vec_tst is
end View_output_vlg_vec_tst;
