library verilog;
use verilog.vl_types.all;
entity Bcd2digitAdder_vlg_vec_tst is
end Bcd2digitAdder_vlg_vec_tst;
