library verilog;
use verilog.vl_types.all;
entity Threebit_BCD_counter_vlg_vec_tst is
end Threebit_BCD_counter_vlg_vec_tst;
