library verilog;
use verilog.vl_types.all;
entity Input_Display_vlg_vec_tst is
end Input_Display_vlg_vec_tst;
