library verilog;
use verilog.vl_types.all;
entity cyclic_reg_with_clock_vlg_vec_tst is
end cyclic_reg_with_clock_vlg_vec_tst;
