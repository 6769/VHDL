library verilog;
use verilog.vl_types.all;
entity adjustAdder4_vlg_vec_tst is
end adjustAdder4_vlg_vec_tst;
