library verilog;
use verilog.vl_types.all;
entity FSM_core_vlg_vec_tst is
end FSM_core_vlg_vec_tst;
