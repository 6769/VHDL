library verilog;
use verilog.vl_types.all;
entity Roll_Sum_vlg_vec_tst is
end Roll_Sum_vlg_vec_tst;
