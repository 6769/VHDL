library verilog;
use verilog.vl_types.all;
entity Counter16anDisplay_vlg_vec_tst is
end Counter16anDisplay_vlg_vec_tst;
