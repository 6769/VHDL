library verilog;
use verilog.vl_types.all;
entity clock_second_vlg_vec_tst is
end clock_second_vlg_vec_tst;
