library verilog;
use verilog.vl_types.all;
entity NumberAnDisplay_vlg_vec_tst is
end NumberAnDisplay_vlg_vec_tst;
